library verilog;
use verilog.vl_types.all;
entity transkoder_vlg_vec_tst is
end transkoder_vlg_vec_tst;
