library verilog;
use verilog.vl_types.all;
entity zad_6_vlg_vec_tst is
end zad_6_vlg_vec_tst;
