library verilog;
use verilog.vl_types.all;
entity zad6_vlg_vec_tst is
end zad6_vlg_vec_tst;
