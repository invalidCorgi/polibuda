library verilog;
use verilog.vl_types.all;
entity skracanie_licznikow_vlg_vec_tst is
end skracanie_licznikow_vlg_vec_tst;
