library verilog;
use verilog.vl_types.all;
entity zad5dudi_vlg_vec_tst is
end zad5dudi_vlg_vec_tst;
